module test_192(
input [191:0] in,
input [31:0] rcon,
output [191:0]out

);
key_expansion_192 key (.key_input(in),.rcon(rcon),.key_output(out));

endmodule 